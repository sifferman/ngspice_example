.lib "$PDK_ROOT/sky130A/libs.tech/combined/sky130.lib.spice" tt
.nodeset all=2.5
.model omod ltra r=1k l=3.333u c=3.333p len=0.02
+ NOCONTROL LININTERP TRUNCNR

VVGND VGND 0 0
VVNB VNB 0 0
VVPB VPB 0 5.0
VVPWR VPWR 0 5.0

.model digital_stimulus d_source(input_file="sky130_fd_sc_hd__dfxtp_1.stim")
a1 [CLK_DIGITAL D_DIGITAL] digital_stimulus

.model dac_model dac_bridge(out_low=0 out_high=5.0 t_rise=2e-11 t_fall=2e-11)
a_dac_bridge1 [CLK_DIGITAL] [CLK] dac_model
a_dac_bridge2 [D_DIGITAL] [D] dac_model

X1 CLK D VGND VNB VPB VPWR Q sky130_fd_sc_hd__dfxtp_1

.control
    tran 10ns 1.2e-06
    wrdata ports.txt CLK D VGND VNB VPB VPWR Q
    exit
.endc

.end
